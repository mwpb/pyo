BZh91AY&SY�G� '߀Px��g߰?���P�䩲��)���x�LmQ�)�'�� �4=A�&0a0�` 2i�a)����SA����z@   �` &	�  &�D� ��O%=G����M�d=OS��=E`b঒��Iy��Iz���f2c�� �C���	 �շ�c��!(��冋D=!�����HEo�H�����XdL"0>�\�:BT��bF��nƖ�ц��鍧����*�}Ή0����a�k��cL�bT
#ͯ��O��:id��x+)�l��"�$щy+&�:�pP�B����&RIb�n�S&Ƭ���a��b4Z�G&�����K�u�}8�
���ƺ��(�.U�;�&�bI#7����z_)밾K꤆��<�Y��������Qj���2�|����B�+��d������xw-<�s#.���B%�k��6��:΀Ρ0m0:e�@�����֦:D��b�����V��|c��ltuhV$!��0`h��3��L�\��ӊ�F�#�D�Cq��KZ�f��T�6���!��\U���c��n��:Y^��;z@�/Z�k�z��KL�@� �u�ު�Y����9q��Y�]��Y�LO	N�9}� �C�2aŽÛ�b1LH�`g  k�цe�j,!P��)�ԗ�a)Z����@��{H=�e�y#�>�����LYvCxV�x�U�5�������-�t�����}����,��p�q�R�.0D�$�7�3lv�܎��/�l�V�o&�'M�i�9K�yl����"�j	�B7^��rN�fr`9dZj��xt�C��L����v0����#�8$WZ��H�
�� 